module main (input  I1, input  I2, input  I3, input  I4, output  D4, output  D3, output  D2, output  D1);
assign D4 = I4;
assign D3 = I3;
assign D2 = I2;
assign D1 = I1;
endmodule

