module main (input [7:0] J1, output [7:0] J3);
wire  inst0_O;
wire  inst1_O;
wire  inst2_O;
wire  inst3_O;
wire  inst4_O;
wire  inst5_O;
wire  inst6_O;
wire  inst7_O;
wire  inst8_O;
wire  inst9_O;
wire  inst10_O;
wire  inst11_O;
wire  inst12_O;
wire  inst13_O;
SB_LUT4 #(.LUT_INIT(16'h9696)) inst0 (.I0(J1[0]), .I1(J1[1]), .I2(J1[2]), .I3(1'b0), .O(inst0_O));
SB_LUT4 #(.LUT_INIT(16'hE8E8)) inst1 (.I0(J1[0]), .I1(J1[1]), .I2(J1[2]), .I3(1'b0), .O(inst1_O));
SB_LUT4 #(.LUT_INIT(16'h9696)) inst2 (.I0(J1[3]), .I1(J1[4]), .I2(J1[5]), .I3(1'b0), .O(inst2_O));
SB_LUT4 #(.LUT_INIT(16'hE8E8)) inst3 (.I0(J1[3]), .I1(J1[4]), .I2(J1[5]), .I3(1'b0), .O(inst3_O));
SB_LUT4 #(.LUT_INIT(16'h9696)) inst4 (.I0(J1[6]), .I1(J1[7]), .I2(1'b0), .I3(1'b0), .O(inst4_O));
SB_LUT4 #(.LUT_INIT(16'hE8E8)) inst5 (.I0(J1[6]), .I1(J1[7]), .I2(1'b0), .I3(1'b0), .O(inst5_O));
SB_LUT4 #(.LUT_INIT(16'h9696)) inst6 (.I0(inst0_O), .I1(inst2_O), .I2(inst4_O), .I3(1'b0), .O(inst6_O));
SB_LUT4 #(.LUT_INIT(16'hE8E8)) inst7 (.I0(inst0_O), .I1(inst2_O), .I2(inst4_O), .I3(1'b0), .O(inst7_O));
SB_LUT4 #(.LUT_INIT(16'h9696)) inst8 (.I0(inst1_O), .I1(inst3_O), .I2(inst5_O), .I3(1'b0), .O(inst8_O));
SB_LUT4 #(.LUT_INIT(16'hE8E8)) inst9 (.I0(inst1_O), .I1(inst3_O), .I2(inst5_O), .I3(1'b0), .O(inst9_O));
SB_LUT4 #(.LUT_INIT(16'h9696)) inst10 (.I0(inst7_O), .I1(inst8_O), .I2(1'b0), .I3(1'b0), .O(inst10_O));
SB_LUT4 #(.LUT_INIT(16'hE8E8)) inst11 (.I0(inst7_O), .I1(inst8_O), .I2(1'b0), .I3(1'b0), .O(inst11_O));
SB_LUT4 #(.LUT_INIT(16'h9696)) inst12 (.I0(inst9_O), .I1(inst10_O), .I2(1'b0), .I3(1'b0), .O(inst12_O));
SB_LUT4 #(.LUT_INIT(16'hE8E8)) inst13 (.I0(inst9_O), .I1(inst10_O), .I2(1'b0), .I3(1'b0), .O(inst13_O));
endmodule

