module main (output  D2, output  D1);
assign D2 = 1'b1;
assign D1 = 1'b1;
endmodule

